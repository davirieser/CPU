
library work;
    use work.CPU_pkg.all;

library ieee;
    use ieee.std_logic_1164.all;


entity Ram is
  port (
    clock   : in std_logic
  );
end Ram;

architecture behaviour of Ram is

    begin

end behaviour;
