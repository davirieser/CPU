library ieee;
	use ieee.std_logic_1164.all;

entity tb_Adder is
end tb_Adder;

architecture behaviour of tb_Adder is

    begin

end behaviour;
