
library work;
    use work.CPU_pkg.all;

library ieee;
    use ieee.std_logic_1164.all;


entity MemoryManager is
  port (
    clock   : in std_logic
  );
end MemoryManager;

architecture behaviour of MemoryManager is

    begin

end behaviour;
