
library work;
    use work.CPU_pkg.all;

library ieee;
    use ieee.std_logic_1164.all;


entity EEPROM is
  port (
    clock   : in std_logic
  );
end EEPROM;

architecture behaviour of EEPROM is

    begin

end behaviour;
