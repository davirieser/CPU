library     ieee;
	use 	ieee.std_logic_1164.all;
	use 	ieee.numeric_std.all;
	use 	ieee.math_real.all;

use work.CPU_pkg.all;

package INST_DEC_pkg is

    -- constant ADD_INST   : std_logic_vector()

end package INST_DEC_pkg;

package body INST_DEC_pkg is

end package body INST_DEC_pkg;
