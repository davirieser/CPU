library work;
    use work.INST_DEC_pkg.all;
    use work.CPU_pkg.all;

library ieee;
	use ieee.std_logic_1164.all;
	use ieee.numeric_std.all;

entity tb_INST_DEC is
end tb_INST_DEC;

architecture behaviour of tb_INST_DEC is

    component INST_DEC is
        port(
            clk         : in std_logic;
            inst        : in std_logic_vector(OPCODE_BITS - 1 downto 0);
            micro_cyc   : in std_logic_vector(NUM_MICRO_CYC - 1 downto 0);
            ctrl_bus    : inout std_logic_vector(ctrl_bus_width - 1 downto 0)
        );
    end component INST_DEC;

    -- 1 + .. => For Clock
    constant size : integer := 1 + OPCODE_BITS + NUM_MICRO_CYC;

    signal sTemp 		: std_logic_vector(size - 1 downto 0) := (others => '0');
    signal sCtrl        : std_logic_vector(ctrl_bus_width - 1 downto 0);

    begin

        uut : entity work.INST_DEC port map(
                                    clk         => sTemp(NUM_MICRO_CYC),
                                    inst        => sTemp(size - 1 downto size - OPCODE_BITS),
                                    micro_cyc   => sTemp(NUM_MICRO_CYC - 1 downto 0),
                                    ctrl_bus    => sCtrl
                                );

		Signal_gen : process

			begin

                for sCount in 0 to (2 ** size) loop

					sTemp <= std_logic_vector(unsigned(sTemp) + 1);

                    wait for base_clock;

                end loop;

				wait;

		end process Signal_gen;

end behaviour;
